module modclk(input wire clk,reset, up, down, output reg z); //z matches modified clock
reg[3:0]state;
parameter A=4'd0,B=4'd1,C=4'd2,D=4'd3,E=4'd4,F=4'd5,G=4'd6,H=4'd7,
I=4'd8,J=4'd9,K=4'd10,L=4'd11;

reg[3:0]next_state;

reg[1/*17*/:0] counter0;//A 0.005s 18bit
reg[2/*18*/:0] counter1;//B 0.01s 19bit
reg[3/*19*/:0] counter2;//C 0.02s 20bit
reg[4/*20*/:0] counter3;//D 0.04s 21bit
reg[5/*21*/:0] counter4;//E 0.08s 22bit
reg[6/*22*/:0] counter5;//F 0.17s 23bit
reg[7/*23*/:0] counter6;//G 0.33s 24bit
reg[8/*24*/:0] counter7;//H 0.67s 25bit
reg[9/*25*/:0] counter8;//I 1.34s 26bit
reg[10/*26*/:0] counter9;//J 2.68s 27bit
reg[11/*27*/:0] counter10;//K 5.36s 28bit
reg[12/*28*/:0] counter11;//L 10.7s 29bit
//12 stats

always @(posedge clk)
if(reset) counter0<=2/*18*/'b0;
else counter0<=counter0+2/*18*/'b1; //~|counter0

always @(posedge clk)
if(reset) counter1<=3/*19*/'b0;
else counter1<=counter1+3/*19*/'b1;

always @(posedge clk)
if(reset) counter2<=4'b0;
else counter2<=counter2+4'b1;

always @(posedge clk)
if(reset) counter3<=5'b0;
else counter3<=counter3+5'b1;

always @(posedge clk)
if(reset) counter4<=6'b0;
else counter4<=counter4+6'b1;
always @(posedge clk)
if(reset) counter5<=7'b0;
else counter5<=counter5+7'b1;

always @(posedge clk)
if(reset) counter6<=24'b0;
else counter6<=counter6+24'b1;

always @(posedge clk)
if(reset) counter7<=8'b0;
else counter7<=counter7+8'b1;

always @(posedge clk)
if(reset) counter8<=9'b0;
else counter8<=counter8+9'b1;

always @(posedge clk)
if(reset) counter9<=10'b0;
else counter9<=counter9+10'b1;

always @(posedge clk)
if(reset) counter10<=11'b0;
else counter10<=counter10+11'b1;

always @(posedge clk)
if(reset) counter11<=12'b0;
else counter11<=counter11+12'b1;

always@(posedge clk)
if(~reset) state<=G;
else state<=next_state;

always@*
case({state,up,down})
{A,1'b1,1'b0}:{next_state,z}={A,~|counter0}; //speed down
{A,1'b0,1'b1}:{next_state,z}={B,~|counter0}; //speed up
{A,1'b0,1'b0}:{next_state,z}={A,~|counter0};
{A,1'b1,1'b1}:{next_state,z}={A,~|counter0};

{B,1'b1,1'b0}:{next_state,z}={A,~|counter1}; //speed down
{B,1'b0,1'b1}:{next_state,z}={C,~|counter1}; //speed up
{B,1'b0,1'b0}:{next_state,z}={B,~|counter1};
{B,1'b1,1'b1}:{next_state,z}={B,~|counter1};

{C,1'b1,1'b0}:{next_state,z}={B,~|counter2}; //speed down
{C,1'b0,1'b1}:{next_state,z}={D,~|counter2}; //speed up
{C,1'b0,1'b0}:{next_state,z}={C,~|counter2};
{C,1'b1,1'b1}:{next_state,z}={C,~|counter2};

{D,1'b1,1'b0}:{next_state,z}={C,~|counter3}; //speed down
{D,1'b0,1'b1}:{next_state,z}={E,~|counter3}; //speed up
{D,1'b0,1'b0}:{next_state,z}={D,~|counter3};
{D,1'b1,1'b1}:{next_state,z}={D,~|counter3};

{E,1'b1,1'b0}:{next_state,z}={D,~|counter4}; //speed down
{E,1'b0,1'b1}:{next_state,z}={F,~|counter4}; //speed up
{E,1'b0,1'b0}:{next_state,z}={E,~|counter4};
{E,1'b1,1'b1}:{next_state,z}={E,~|counter4};

{F,1'b1,1'b0}:{next_state,z}={E,~|counter5}; //speed down
{F,1'b0,1'b1}:{next_state,z}={G,~|counter5}; //speed up
{F,1'b0,1'b0}:{next_state,z}={F,~|counter5};
{F,1'b1,1'b1}:{next_state,z}={F,~|counter5};

{G,1'b1,1'b0}:{next_state,z}={F,~|counter6}; //speed down
{G,1'b0,1'b1}:{next_state,z}={H,~|counter6}; //speed up
{G,1'b0,1'b0}:{next_state,z}={G,~|counter6};
{G,1'b1,1'b1}:{next_state,z}={G,~|counter6};

{H,1'b1,1'b0}:{next_state,z}={G,~|counter7}; //speed down
{H,1'b0,1'b1}:{next_state,z}={I,~|counter7}; //speed up
{H,1'b0,1'b0}:{next_state,z}={H,~|counter7};
{H,1'b1,1'b1}:{next_state,z}={H,~|counter7};

{I,1'b1,1'b0}:{next_state,z}={H,~|counter8}; //speed down
{I,1'b0,1'b1}:{next_state,z}={J,~|counter8}; //speed up
{I,1'b0,1'b0}:{next_state,z}={I,~|counter8};
{I,1'b1,1'b1}:{next_state,z}={I,~|counter8};

{J,1'b1,1'b0}:{next_state,z}={I,~|counter9}; //speed down
{J,1'b0,1'b1}:{next_state,z}={K,~|counter9}; //speed up
{J,1'b0,1'b0}:{next_state,z}={J,~|counter9};
{J,1'b1,1'b1}:{next_state,z}={J,~|counter9};

{K,1'b1,1'b0}:{next_state,z}={J,~|counter10}; //speed down
{K,1'b0,1'b1}:{next_state,z}={L,~|counter10}; //speed up
{K,1'b0,1'b0}:{next_state,z}={K,~|counter10};
{K,1'b1,1'b1}:{next_state,z}={K,~|counter10};

{L,1'b1,1'b0}:{next_state,z}={K,~|counter11}; //speed down
{L,1'b0,1'b1}:{next_state,z}={L,~|counter11}; //speed up
{L,1'b0,1'b0}:{next_state,z}={L,~|counter11};
{L,1'b1,1'b1}:{next_state,z}={L,~|counter11};
default:{next_state,z}={G,~|counter6};     //Default goes to G state (0.33s)
endcase
endmodule
