module DEC13(input wire[6:0]i,output reg[6:0]o);
always @*
case(i)
7'd0: o=7'b1111111;
7'd1: o=7'b1111111;
7'd2: o=7'b1111111;
7'd3: o=7'b1111111;
7'd4: o=7'b1111111;
7'd5: o=7'b1110111;
7'd6: o=7'b1110111;
7'd7: o=7'b1110111;
7'd8: o=7'b1111111;
7'd9: o=7'b1111111;
7'd10:o=7'b1111111;
7'd11:o=7'b1111111;
7'd12:o=7'b1111111;
7'd13:o=7'b1111111;
7'd14:o=7'b1111111;
7'd15:o=7'b1111111;
7'd16:o=7'b1111111;
7'd17:o=7'b1111111;
7'd18:o=7'b1111111;
7'd19:o=7'b1111111;
7'd20:o=7'b1111111;
7'd21:o=7'b1011111;
7'd22:o=7'b1011101;
7'd23:o=7'b1011111;
7'd24:o=7'b1111111;
7'd25:o=7'b1111111;
7'd26:o=7'b1111111;
7'd27:o=7'b1111111;
7'd28:o=7'b1111111;
7'd29:o=7'b1111111;
7'd30:o=7'b1111111;
7'd31:o=7'b1111111;
7'd32:o=7'b1111111;
7'd33:o=7'b1111111;
7'd34:o=7'b1111111;
7'd35:o=7'b1111111;
7'd36:o=7'b1111111;
7'd37:o=7'b1111110;
7'd38:o=7'b1111111;
7'd39:o=7'b1111111;
7'd40:o=7'b1111111;
7'd41:o=7'b1111111;
7'd42:o=7'b1111111;
7'd43:o=7'b1111111;
7'd44:o=7'b1111111;
7'd45:o=7'b1111111;
7'd46:o=7'b1111111;
7'd47:o=7'b1111111;
7'd48:o=7'b1111111;
7'd49:o=7'b1111111;
7'd50:o=7'b1111111;
7'd51:o=7'b1101111;
7'd52:o=7'b1101011;
7'd53:o=7'b1101011;
7'd54:o=7'b1101011;
7'd55:o=7'b1101111;
7'd56:o=7'b1111111;
7'd57:o=7'b1111111;
7'd58:o=7'b1111111;
7'd59:o=7'b1111111;
7'd60:o=7'b1111111;
7'd61:o=7'b1111111;
7'd62:o=7'b1111111;
7'd63:o=7'b1111111;
7'd64:o=7'b1111111;
7'd65:o=7'b1111111;
7'd66:o=7'b1111111;
7'd67:o=7'b1111111;
7'd68:o=7'b1111111;
7'd69:o=7'b0111111;
7'd70:o=7'b0111111;
7'd71:o=7'b0111111;
7'd72:o=7'b1111111;
7'd73:o=7'b1111111;
7'd74:o=7'b1111111;
7'd75:o=7'b1111111;
7'd76:o=7'b1111111;
7'd77:o=7'b1111111;
7'd78:o=7'b1111111;
7'd79:o=7'b1111111;
7'd80:o=7'b1111111;
7'd81:o=7'b1111111;
7'd82:o=7'b1111111;
7'd83:o=7'b1111111;
7'd84:o=7'b1111111;
7'd85:o=7'b1111111;
7'd86:o=7'b1111111;
7'd87:o=7'b1111111;
7'd88:o=7'b1111111;
7'd89:o=7'b1111111;
7'd90:o=7'b1111111;
7'd91:o=7'b1111111;
7'd92:o=7'b1111111;
7'd93:o=7'b1111111;
7'd94:o=7'b1111111;
7'd95:o=7'b1111111;
7'd96:o=7'b1111111;
7'd97:o=7'b0110110;
7'd98:o=7'b0110110;
7'd99:o=7'b0110110;
7'd100:o=7'b1111111;
7'd101:o=7'b1111111;
7'd102:o=7'b1111111;
7'd103:o=7'b1111111;
7'd104:o=7'b1111111;
7'd105:o=7'b1111111;
7'd106:o=7'b1111111;
7'd107:o=7'b1111111;
7'd108:o=7'b1111111;
7'd109:o=7'b1111111;
7'd110:o=7'b1111111;
7'd111:o=7'b1111111;
7'd112:o=7'b1111111;
7'd113:o=7'b1001111;
7'd114:o=7'b1001001;
7'd115:o=7'b1001001;
7'd116:o=7'b1001001;
7'd117:o=7'b1001001;
7'd118:o=7'b1001001;
7'd119:o=7'b1001111;
7'd120:o=7'b1111111;
7'd121:o=7'b1111111;
7'd122:o=7'b1111111;
7'd123:o=7'b1111111;
7'd124:o=7'b1111111;
7'd125:o=7'b1111111;
7'd126:o=7'b1111111;
7'd127:o=7'b1111111;
endcase 
endmodule
