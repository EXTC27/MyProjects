module LED_DEC0(input wire[4:0]i,output reg[9:0]o);
always @*
case(i)
5'd0: o=10'b0000000000;//0 meas out 1 means bright
5'd1: o=10'b1000000000;
5'd2: o=10'b1100000000;
5'd3: o=10'b1110000000;
5'd4: o=10'b1111000000;
5'd5: o=10'b1111100000;
5'd6: o=10'b1111110000;
5'd7: o=10'b1111111000;
5'd8: o=10'b1111111100;
5'd9: o=10'b1111111110;
5'd10:o=10'b1111111111;
5'd11:o=10'b1111111110;
5'd12:o=10'b1111111100;
5'd13:o=10'b1111111000;
5'd14:o=10'b1111110000;
5'd15:o=10'b1111100000;
5'd16:o=10'b1111000000;
5'd17:o=10'b1110000000;
5'd18:o=10'b1100000000;
5'd19:o=10'b1000000000;
5'd20:o=10'b0000000000;
5'd21:o=10'b1000000000;
5'd22:o=10'b1100000000;
5'd23:o=10'b1110000000;
5'd24:o=10'b1111000000;
5'd25:o=10'b1111100000;
5'd26:o=10'b1111000000;
5'd27:o=10'b1110000000;
5'd28:o=10'b1100000000;
5'd29:o=10'b1000000000;
5'd30:o=10'b0000000000;
5'd31:o=10'b0000000000;
endcase 
endmodule
